
 
 module truckBitMap (

					input	logic	clk, 
					input	logic	resetN, 
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY, 
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
 
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ; 
 
 
// generating the bitmap 
 

localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel  
logic[0:63][127:0][7:0] object_colors = {
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'hfb,8'hfb,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'hfb,8'hfb,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'hfb,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'hd7,8'h00,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hdf,8'hbb,8'h97,8'h77,8'h97,8'h32,8'h72,8'h32,8'h2e,8'h32,8'h72,8'h32,8'h73,8'h32,8'h32,8'h33,8'h32,8'h37,8'h32,8'h32,8'h37,8'h32,8'h32,8'h32,8'h2e,8'h97,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hbb,8'h73,8'h72,8'h2e,8'h2e,8'h2e,8'h2e,8'h2e,8'h2e,8'h2e,8'h2e,8'h2e,8'h2e,8'h2e,8'h2e,8'h2e,8'h2e,8'h72,8'h73,8'h93,8'hb7,8'hbb,8'hdb,8'hdf,8'h00,8'h00,8'h00,8'hfb,8'hfb,8'hd7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'hd7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h73,8'h2e,8'h0e,8'h32,8'h77,8'h32,8'h12,8'h32,8'h33,8'h77,8'h77,8'h32,8'h77,8'h77,8'h33,8'h77,8'h33,8'h33,8'h37,8'h33,8'h77,8'h37,8'h37,8'h77,8'h37,8'h37,8'h37,8'h32,8'h32,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h73,8'h2e,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h2e,8'h2e,8'h2e,8'h32,8'h2e,8'h2e,8'h72,8'h93,8'hb7,8'hdb,8'h00,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h77,8'h37,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h37,8'h77,8'h7b,8'h7b,8'h9b,8'h9b,8'hbb,8'hbb,8'h9b,8'hbb,8'hbb,8'h9b,8'h9b,8'h77,8'h7b,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h37,8'h37,8'h33,8'h32,8'h32,8'h32,8'h73,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h73,8'h2e,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h0e,8'h32,8'h32,8'h0e,8'hbb,8'h77,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h12,8'h12,8'h12,8'h32,8'h32,8'h37,8'h37,8'h37,8'h77,8'h77,8'h77,8'h7b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h77,8'h77,8'h77,8'h33,8'h33,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h93,8'hdb,8'h00,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hd7,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h77,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h77,8'hbf,8'hbf,8'hbf,8'hbf,8'hbf,8'hbb,8'hbb,8'hbf,8'hbb,8'hbb,8'hbb,8'hbb,8'hbf,8'hbf,8'hbb,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h32,8'h12,8'h37,8'h37,8'h32,8'h37,8'h33,8'h37,8'h37,8'h32,8'h37,8'h37,8'h37,8'h77,8'h33,8'h77,8'h37,8'h32,8'h32,8'h32,8'h32,8'h73,8'h77,8'h33,8'h32,8'h32,8'h32,8'h32,8'h32,8'h33,8'h37,8'h37,8'h37,8'h77,8'h77,8'h32,8'h77,8'h37,8'h37,8'h37,8'h32,8'h32,8'h12,8'h32,8'h37,8'h37,8'h37,8'h37,8'h37,8'h9f,8'hbf,8'hbf,8'hbf,8'hbf,8'hbf,8'hbf,8'hbf,8'hbf,8'hbf,8'hbf,8'hbf,8'hbf,8'hbf,8'hbf,8'hbb,8'hbb,8'h9b,8'h9b,8'h77,8'h37,8'h33,8'h32,8'h32,8'h77,8'hbb,8'hdb,8'hb3,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hd7,8'h00,8'hfb,8'hfb,8'h00,8'h00,8'hbb,8'h37,8'h37,8'h37,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h33,8'h33,8'h32,8'h33,8'h33,8'h37,8'h37,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h12,8'h32,8'h33,8'h32,8'h12,8'h32,8'h32,8'h72,8'h72,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h33,8'h33,8'h33,8'h37,8'h33,8'h33,8'h77,8'h37,8'h37,8'h37,8'h37,8'h32,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h33,8'h33,8'h33,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h7b,8'h37,8'h77,8'hdb,8'h72,8'hdb,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hd7,8'hfb,8'hfb,8'h93,8'h00,8'h00,8'h97,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h33,8'h33,8'h0d,8'h0e,8'h37,8'h37,8'h32,8'h2e,8'h0e,8'h2e,8'h2e,8'h2e,8'h2e,8'h32,8'h2e,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h9b,8'h9b,8'h32,8'h32,8'h32,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h37,8'h37,8'h37,8'h73,8'hbb,8'h32,8'h00,8'hd7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb3,8'hfb,8'h92,8'hb7,8'h97,8'h97,8'h97,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h9b,8'h77,8'h9b,8'h37,8'h32,8'h33,8'h37,8'h37,8'h37,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h33,8'h77,8'h33,8'h32,8'h32,8'h37,8'h37,8'h12,8'h12,8'h12,8'h12,8'h13,8'h12,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h73,8'h77,8'h77,8'h00,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'hfb,8'hb7,8'h9b,8'h77,8'h9b,8'h7b,8'h7b,8'h9b,8'h7b,8'h9b,8'h9b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h9b,8'h77,8'h9b,8'h33,8'h32,8'h37,8'h37,8'h37,8'h37,8'h77,8'h37,8'h37,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h33,8'h37,8'h37,8'h33,8'h77,8'h77,8'h0e,8'h0d,8'h0d,8'h2e,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h17,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h33,8'h73,8'h00,8'hd7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hd7,8'hfb,8'h00,8'h97,8'h32,8'h37,8'h37,8'h32,8'h37,8'h33,8'h32,8'h33,8'h33,8'h33,8'h37,8'h37,8'h32,8'h33,8'h37,8'h37,8'h37,8'h33,8'h33,8'h32,8'h32,8'h33,8'h33,8'h33,8'h37,8'h37,8'h33,8'h33,8'h37,8'h37,8'h33,8'h33,8'h33,8'h33,8'h33,8'h37,8'h37,8'h33,8'h37,8'h37,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h33,8'h9b,8'h33,8'h32,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h77,8'h77,8'h77,8'h77,8'h77,8'h7b,8'h7b,8'h7b,8'h77,8'h33,8'h37,8'h32,8'h0d,8'h25,8'h2e,8'h2e,8'h32,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h17,8'h16,8'h12,8'h12,8'h16,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h77,8'h37,8'hbb,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb3,8'hfb,8'h00,8'h97,8'h12,8'h37,8'h12,8'h37,8'h17,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h33,8'h37,8'h32,8'h33,8'h32,8'h32,8'h33,8'h32,8'h9b,8'h77,8'h32,8'h37,8'h17,8'h37,8'h37,8'h7b,8'h3b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h77,8'h37,8'h32,8'h05,8'h25,8'h6e,8'h2e,8'h32,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h17,8'h12,8'h12,8'h17,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h12,8'h9b,8'h37,8'h33,8'h97,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hd7,8'hfb,8'h00,8'h97,8'h37,8'h17,8'h33,8'h37,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h32,8'h32,8'h32,8'h9b,8'h77,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h77,8'h77,8'h77,8'h77,8'h77,8'h77,8'h7b,8'h7b,8'h7b,8'h37,8'h73,8'h05,8'h25,8'h65,8'h2e,8'h32,8'h32,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h13,8'h12,8'h12,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h12,8'hbb,8'h37,8'h37,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hd7,8'hfb,8'h00,8'h97,8'h36,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h32,8'h32,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h77,8'h0d,8'h25,8'h25,8'h6e,8'h2e,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h12,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h33,8'h12,8'hbf,8'h37,8'h37,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hd7,8'hfb,8'h00,8'h97,8'h33,8'h12,8'h33,8'h37,8'h17,8'h17,8'h37,8'h37,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h32,8'h32,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h77,8'h2e,8'h25,8'h25,8'h6e,8'h32,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h7b,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h12,8'h12,8'h37,8'h33,8'h37,8'h37,8'h12,8'hbf,8'h37,8'h37,8'h32,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'hb7,8'h97,8'h37,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h32,8'h32,8'h7b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h9b,8'h73,8'h32,8'h25,8'h25,8'h2e,8'h2d,8'h37,8'h37,8'h37,8'h37,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h7b,8'h7b,8'h7b,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h32,8'h32,8'h32,8'h12,8'hbf,8'h37,8'h37,8'h73,8'hbb,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb3,8'hfb,8'h97,8'h77,8'h32,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h32,8'h32,8'h7b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h73,8'h72,8'h25,8'h25,8'h6e,8'h05,8'h33,8'h37,8'h37,8'h37,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h7b,8'h7b,8'h7b,8'h77,8'h37,8'h37,8'h37,8'h37,8'h12,8'h32,8'h32,8'h12,8'h0e,8'hbf,8'h33,8'h37,8'h73,8'hb7,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h32,8'h17,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h32,8'h32,8'h7b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h77,8'h72,8'h25,8'h25,8'h6e,8'h25,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h77,8'h7b,8'h9b,8'h7b,8'h37,8'h37,8'h37,8'h37,8'h12,8'h32,8'h33,8'h33,8'h37,8'h37,8'h33,8'h97,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h12,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h37,8'h37,8'h37,8'h37,8'h37,8'h32,8'h32,8'h7b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h77,8'h73,8'h25,8'h25,8'h6e,8'h25,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h7b,8'h37,8'h37,8'h37,8'h12,8'h12,8'h33,8'h32,8'h9b,8'h37,8'h33,8'h97,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h12,8'h17,8'h37,8'h37,8'h37,8'h37,8'h17,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h77,8'h73,8'h25,8'h25,8'h6e,8'h25,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h77,8'h37,8'h33,8'h32,8'h32,8'h32,8'h9b,8'h9b,8'h33,8'h77,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h12,8'h13,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h77,8'h73,8'h25,8'h25,8'h2e,8'h2d,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h7b,8'h37,8'h32,8'h32,8'h32,8'h32,8'h33,8'hbf,8'h77,8'h73,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h33,8'h12,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h77,8'h77,8'h25,8'h25,8'h6e,8'h2e,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h37,8'h37,8'h7b,8'h7b,8'h7b,8'h7b,8'h37,8'h33,8'h12,8'h32,8'h12,8'h7b,8'h73,8'h73,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h32,8'h13,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h77,8'h77,8'h25,8'h25,8'h6e,8'h6e,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h37,8'h37,8'h9b,8'h7b,8'h9b,8'h9b,8'h37,8'h37,8'h12,8'h12,8'h12,8'h77,8'h32,8'h73,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h37,8'h12,8'h37,8'h37,8'h37,8'h17,8'h12,8'h17,8'h17,8'h17,8'h37,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h77,8'h77,8'h25,8'h25,8'h2e,8'h6e,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h37,8'h37,8'h37,8'h9b,8'h7b,8'h9b,8'h77,8'h37,8'h37,8'h12,8'h12,8'h32,8'h32,8'h32,8'h73,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h33,8'h13,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h77,8'h77,8'h25,8'h25,8'h6e,8'h6e,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h37,8'h37,8'h37,8'h7b,8'h77,8'h9b,8'h77,8'h37,8'h37,8'h12,8'h12,8'h12,8'h32,8'h77,8'h73,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h33,8'h13,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h77,8'h77,8'h25,8'h25,8'h6e,8'h6e,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h9b,8'h97,8'h77,8'h77,8'h37,8'h12,8'h12,8'h12,8'h32,8'h97,8'h72,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h32,8'h13,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h77,8'h77,8'h25,8'h25,8'h6e,8'h6e,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h9b,8'h97,8'h9b,8'h7b,8'h37,8'h12,8'h16,8'h32,8'h12,8'h97,8'h73,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h32,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h77,8'h77,8'h25,8'h25,8'h6e,8'h6e,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h9b,8'h77,8'h9b,8'h7b,8'h37,8'h12,8'h16,8'h32,8'h32,8'h97,8'h72,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h32,8'h13,8'h37,8'h37,8'h37,8'h37,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h77,8'h77,8'h25,8'h25,8'h6e,8'h6e,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h97,8'h9b,8'h77,8'h37,8'h12,8'h16,8'h12,8'h12,8'h97,8'h73,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h33,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h77,8'h77,8'h25,8'h25,8'h6e,8'h6e,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h9b,8'h77,8'h9b,8'h77,8'h37,8'h37,8'h12,8'h12,8'h32,8'h12,8'h73,8'h73,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h33,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h32,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h77,8'h77,8'h25,8'h25,8'h6e,8'h6e,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h9b,8'h77,8'h33,8'h37,8'h12,8'h12,8'h32,8'h32,8'h32,8'h73,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h33,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h77,8'h77,8'h25,8'h25,8'h6e,8'h6e,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h7b,8'h7b,8'h37,8'h37,8'h12,8'h32,8'h12,8'h77,8'h73,8'h73,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hd7,8'hfb,8'h00,8'h97,8'h32,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h77,8'h77,8'h25,8'h25,8'h6e,8'h2d,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h77,8'h37,8'h32,8'h12,8'h12,8'h33,8'h12,8'hbf,8'h77,8'h73,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hd7,8'hfb,8'h00,8'h97,8'h32,8'h12,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h7b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h9b,8'h77,8'h73,8'h25,8'h25,8'h6e,8'h25,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h77,8'h37,8'h37,8'h12,8'h12,8'h32,8'h77,8'h9f,8'h77,8'h73,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h33,8'h12,8'h16,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h7b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h37,8'h37,8'h37,8'h7b,8'h9b,8'h77,8'h73,8'h25,8'h25,8'h6e,8'h25,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h7b,8'h37,8'h37,8'h37,8'h12,8'h12,8'h32,8'h9f,8'h77,8'h33,8'h97,8'hd7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h32,8'h17,8'h12,8'h37,8'h37,8'h37,8'h17,8'h17,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h17,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h77,8'h32,8'h25,8'h25,8'h6e,8'h2d,8'h77,8'h37,8'h37,8'h37,8'h37,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h7b,8'h77,8'h37,8'h37,8'h37,8'h12,8'h32,8'h32,8'h32,8'h7b,8'h37,8'h37,8'h97,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hd7,8'hfb,8'h00,8'h97,8'h32,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h77,8'h77,8'h32,8'h25,8'h25,8'h6e,8'h05,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h7b,8'h7b,8'h77,8'h37,8'h37,8'h37,8'h12,8'h12,8'h32,8'h32,8'h77,8'h37,8'h37,8'h37,8'h97,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h97,8'h97,8'h37,8'h16,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h32,8'h32,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h73,8'h32,8'h25,8'h25,8'h6e,8'h2d,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h7b,8'h7b,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h32,8'h32,8'h12,8'hbf,8'h37,8'h37,8'h33,8'hb7,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'hdf,8'h97,8'h12,8'h37,8'h37,8'h37,8'h37,8'h17,8'h17,8'h17,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h37,8'h37,8'h37,8'h17,8'h17,8'h17,8'h17,8'h37,8'h37,8'h32,8'h32,8'h9b,8'h37,8'h12,8'h37,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h77,8'h2e,8'h25,8'h25,8'h2e,8'h2e,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h7b,8'h7b,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h12,8'h12,8'h32,8'h32,8'h12,8'hbf,8'h37,8'h37,8'h37,8'hbb,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h32,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h32,8'h32,8'h9b,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h77,8'h2e,8'h25,8'h25,8'h6e,8'h2e,8'h37,8'h37,8'h37,8'h37,8'h17,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h7b,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h33,8'h12,8'h12,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'hbf,8'h37,8'h37,8'h32,8'hdf,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h36,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h32,8'h32,8'h9b,8'h77,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h77,8'h77,8'h0d,8'h25,8'h25,8'h6e,8'h2e,8'h12,8'h37,8'h37,8'h17,8'h17,8'h17,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h12,8'h16,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h32,8'h12,8'hbf,8'h37,8'h37,8'h73,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb3,8'hfb,8'h00,8'h97,8'h32,8'h12,8'h12,8'h16,8'h17,8'h17,8'h12,8'h37,8'h12,8'h12,8'h12,8'h17,8'h37,8'h32,8'h12,8'h12,8'h12,8'h16,8'h16,8'h12,8'h12,8'h12,8'h12,8'h12,8'h13,8'h13,8'h12,8'h12,8'h13,8'h33,8'h32,8'h32,8'h32,8'h32,8'h32,8'h33,8'h33,8'h33,8'h32,8'h12,8'h12,8'h12,8'h32,8'h33,8'h32,8'h32,8'h32,8'h97,8'h73,8'h32,8'h37,8'h37,8'h37,8'h37,8'h3b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h37,8'h32,8'h05,8'h25,8'h25,8'h2e,8'h32,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h12,8'h12,8'h16,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h12,8'h12,8'h9b,8'h37,8'h37,8'h97,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h32,8'h32,8'h37,8'h17,8'h17,8'h37,8'h37,8'h37,8'h33,8'h37,8'h37,8'h33,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h33,8'h33,8'h33,8'h33,8'h33,8'h33,8'h33,8'h33,8'h33,8'h33,8'h33,8'h32,8'h9b,8'h77,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h37,8'h37,8'h32,8'h25,8'h25,8'h66,8'h2e,8'h32,8'h37,8'h37,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h12,8'h12,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h12,8'hbf,8'h37,8'h33,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h97,8'h77,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h33,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h37,8'h37,8'h0d,8'h05,8'h25,8'h2e,8'h32,8'h32,8'h37,8'h37,8'h37,8'h37,8'h37,8'h33,8'h32,8'h33,8'h13,8'h12,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h17,8'h17,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h33,8'h97,8'h37,8'h77,8'hdb,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'hb7,8'h97,8'h97,8'h97,8'h97,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h9b,8'h7b,8'h77,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h33,8'h32,8'h33,8'h37,8'h37,8'h37,8'h37,8'h33,8'h73,8'h77,8'h37,8'h77,8'h33,8'h33,8'h73,8'h73,8'h73,8'h73,8'h33,8'h33,8'h73,8'h37,8'h77,8'h32,8'h2e,8'h2d,8'h2e,8'h33,8'h37,8'h37,8'h37,8'h13,8'h13,8'h12,8'h12,8'h12,8'h12,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h33,8'h33,8'h00,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb3,8'hfb,8'h93,8'h97,8'h97,8'h97,8'h97,8'h77,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h77,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h77,8'h77,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h33,8'h32,8'h33,8'h37,8'h37,8'h33,8'h32,8'h2e,8'h2e,8'h2e,8'h0e,8'h0e,8'h0d,8'h0d,8'h0d,8'h0d,8'h0d,8'h0d,8'h0d,8'h0e,8'h0e,8'h32,8'h32,8'h73,8'h73,8'h73,8'h73,8'h37,8'h17,8'h12,8'h12,8'h12,8'h12,8'h13,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h73,8'h97,8'h73,8'h00,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'hb7,8'h00,8'h00,8'hbb,8'h37,8'h37,8'h37,8'h36,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h0e,8'h12,8'h32,8'h33,8'h33,8'h2e,8'h2e,8'h2e,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h33,8'h32,8'h73,8'h9b,8'h77,8'h37,8'h33,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h33,8'h33,8'h37,8'h37,8'h37,8'h37,8'h33,8'h73,8'hdb,8'h72,8'h00,8'hd7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hd7,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'h37,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h7b,8'h77,8'h77,8'h77,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h33,8'h37,8'h37,8'h32,8'h32,8'h12,8'h32,8'h33,8'h77,8'h73,8'h32,8'h32,8'h32,8'h33,8'h33,8'h33,8'h33,8'h33,8'h33,8'h37,8'h37,8'h77,8'h33,8'h33,8'h9b,8'h33,8'h12,8'h37,8'h33,8'h12,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h77,8'h7b,8'h7b,8'h9b,8'h9b,8'h9b,8'h9f,8'h9f,8'h9f,8'h9b,8'h9b,8'h33,8'h97,8'hdb,8'h93,8'hdb,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hfb,8'hd7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h32,8'h32,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h7b,8'h9b,8'h9b,8'hbf,8'hbf,8'hbf,8'hbf,8'hbb,8'hbb,8'hbf,8'hbf,8'hbf,8'hbf,8'h9b,8'h9b,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h32,8'h12,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h33,8'h12,8'h77,8'h32,8'h33,8'h32,8'h33,8'h33,8'h33,8'h32,8'h32,8'h32,8'h33,8'h37,8'h37,8'h33,8'h37,8'h77,8'h9b,8'h9b,8'h9b,8'h9b,8'h9f,8'hbf,8'hbf,8'hbf,8'hbf,8'hbf,8'hbb,8'h9b,8'h9b,8'h9b,8'h77,8'h77,8'h37,8'h33,8'h32,8'h32,8'h32,8'h32,8'h32,8'h93,8'hbb,8'hdb,8'hb7,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb7,8'hd7,8'h00,8'h00,8'h00,8'h00,8'h97,8'h32,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h77,8'h7b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h9b,8'h77,8'h77,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h12,8'h12,8'h32,8'h0e,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h2e,8'h2e,8'h32,8'h32,8'h32,8'h32,8'h2e,8'h2e,8'h32,8'h32,8'h32,8'h32,8'h0d,8'hbb,8'h97,8'h32,8'h0e,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h33,8'h33,8'h33,8'h33,8'h33,8'h33,8'h33,8'h33,8'h33,8'h33,8'h32,8'h32,8'h32,8'h33,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h73,8'hdb,8'h00,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'hbb,8'h97,8'h32,8'h32,8'h32,8'h32,8'h0e,8'h0e,8'h32,8'h32,8'h32,8'h32,8'h33,8'h33,8'h33,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h37,8'h33,8'h32,8'h32,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'h97,8'h2e,8'h2e,8'h2e,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h2e,8'h2e,8'h2e,8'h2e,8'h73,8'h97,8'hbb,8'hbb,8'h00,8'hdb,8'h00,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'hb7,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdf,8'hdb,8'h97,8'h97,8'h73,8'h73,8'h32,8'h0e,8'h2e,8'h2e,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h0e,8'h2e,8'h73,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hbb,8'h97,8'h93,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h73,8'h73,8'h73,8'h97,8'hb7,8'hb7,8'hdb,8'hdb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb3,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hfb,8'h00,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'h00,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}};

 
 

//////////--------------------------------------------------------------------------------------------------------------= 
always_ff@(posedge clk or negedge resetN) 
begin 
	if(!resetN) begin 
		RGBout <=	8'h00; 
	end 
	else begin 
		RGBout <= TRANSPARENT_ENCODING ; // default  
 
		if (InsideRectangle == 1'b1 ) 
		begin // inside an external bracket  
			RGBout <= object_colors[offsetX][offsetY]; 
		end  	 
		 
	end 
end 
 
//////////--------------------------------------------------------------------------------------------------------------= 
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
 
endmodule 
