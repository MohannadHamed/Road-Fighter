
 module introPicBitMap (

					input	logic	clk, 
					input	logic	resetN, 
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY, 
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ; 
 
 
// generating the bitmap 
 

localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel  
logic[0:127][0:127][7:0] object_colors = {
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hda,8'hda,8'hff,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hda,8'hff,8'hda,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hda,8'hff,8'hff,8'hff,8'hda,8'hff,8'hda,8'hda,8'hda,8'hff,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'hb6,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'hb6,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hb6,8'h91,8'h2d,8'h35,8'h35,8'h35,8'h35,8'h36,8'h36,8'h36,8'h36,8'h36,8'h35,8'h36,8'h36,8'h36,8'hd4,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf8,8'h35,8'h2d,8'h35,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h35,8'h35,8'h35,8'h00,8'h8c,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h91,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hb6,8'h31,8'h36,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7e,8'h7a,8'h7e,8'h7e,8'h7a,8'h9a,8'hfc,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h24,8'h24,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h35,8'h35,8'h36,8'h36,8'h35,8'h35,8'h35,8'h35,8'h36,8'h00,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h8c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'h35,8'h7a,8'h7a,8'h7a,8'h7a,8'h9a,8'hf9,8'hfc,8'hfc,8'hd4,8'h24,8'h24,8'h91,8'hda,8'hda,8'hb6,8'h91,8'h91,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd8,8'h35,8'h35,8'h36,8'h36,8'h36,8'h00,8'hfc,8'hfc,8'hfc,8'hf8,8'hfc,8'hf8,8'hfc,8'hfc,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'h7a,8'h7a,8'hfc,8'h00,8'h91,8'hff,8'hff,8'hda,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h6d,8'h00,8'h24,8'h6d,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd8,8'h35,8'h36,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h6d,8'h91,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7a,8'hda,8'hda,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hda,8'h24,8'h00,8'h00,8'h91,8'hb6,8'h91,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h00,8'h00,8'h00,8'h6d,8'h24,8'h91,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h00,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h9a,8'h7a,8'h7a,8'h7a,8'hfc,8'hb6,8'h24,8'hda,8'hb6,8'hb6,8'h00,8'h91,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'h24,8'h24,8'hb6,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'h00,8'h24,8'h6d,8'h6d,8'hb6,8'hb6,8'h91,8'h91,8'h91,8'h91,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h9a,8'h7a,8'h7a,8'h7a,8'h7a,8'h6d,8'h24,8'h91,8'h00,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'h00,8'h00,8'h6d,8'h91,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h91,8'h91,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb0,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdf,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h24,8'h00,8'h91,8'h6d,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'h00,8'h91,8'h6d,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h91,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf8,8'h24,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'hfd,8'h00,8'h24,8'h24,8'h91,8'h24,8'h91,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hff,8'h6d,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfc,8'hb0,8'h91,8'h91,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'hb6,8'h91,8'h91,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h36,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h9a,8'hda,8'hff,8'h24,8'h24,8'h24,8'h6d,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfc,8'h90,8'h91,8'hda,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hf8,8'h00,8'h6d,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h36,8'h35,8'h7a,8'h7a,8'h7a,8'h7e,8'h7e,8'h7e,8'hfc,8'hda,8'hff,8'h91,8'h6d,8'h24,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h24,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfc,8'h6d,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf8,8'hd4,8'h00,8'h24,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h35,8'h35,8'h35,8'h36,8'h7a,8'h7a,8'h7a,8'h7e,8'hd9,8'h24,8'hda,8'h00,8'h6d,8'h24,8'h24,8'h24,8'hff,8'hff,8'hff,8'hb6,8'h6d,8'h6d,8'h6d,8'h24,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'h91,8'h00,8'hfc,8'h6d,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h9a,8'h35,8'h35,8'h35,8'h35,8'h36,8'h36,8'h7e,8'h7e,8'h7a,8'hfc,8'hff,8'hff,8'h00,8'h24,8'h00,8'h00,8'h6d,8'hff,8'h24,8'h91,8'h6d,8'h24,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb0,8'h6d,8'h24,8'h00,8'h00,8'hfc,8'h00,8'h6d,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h91,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00},
	{8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h35,8'h2d,8'h35,8'h35,8'h35,8'h36,8'h36,8'h35,8'h36,8'h7e,8'h7e,8'hfc,8'hda,8'hff,8'h00,8'h00,8'h00,8'h00,8'h91,8'h24,8'h24,8'h6d,8'h6d,8'h24,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'h6d,8'h24,8'h00,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'h6d,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hf8,8'h00,8'h00,8'h91,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00},
	{8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h35,8'h2d,8'h35,8'h35,8'h35,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h7e,8'hd9,8'hb6,8'hff,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h24,8'h24,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h24,8'h00,8'h24,8'h00,8'h00,8'h00,8'h24,8'h00,8'h6d,8'h6d,8'h6d,8'h00,8'h24,8'h00,8'h00,8'hfc,8'hfc,8'h6d,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00},
	{8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h2d,8'h35,8'h35,8'h36,8'h35,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'hfc,8'h00,8'hda,8'hff,8'h00,8'h00,8'h00,8'h00,8'h91,8'h24,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h00,8'h6d,8'h00,8'h00,8'h24,8'h24,8'h00,8'h00,8'hfc,8'h00,8'h6d,8'hb6,8'h91,8'hb6,8'h91,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00},
	{8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h31,8'h2d,8'h35,8'h35,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'hfc,8'h00,8'hda,8'hff,8'h00,8'h00,8'h6d,8'h24,8'h6d,8'h00,8'h24,8'h24,8'h00,8'h24,8'h00,8'h24,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h00,8'h00,8'h8c,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'h00,8'hfc,8'hfc,8'h6d,8'hb6,8'h91,8'h91,8'h91,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'h00,8'hd4,8'hd4,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00},
	{8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h35,8'h35,8'h35,8'h35,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'hfc,8'h24,8'hda,8'hff,8'h00,8'h91,8'h00,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h91,8'h24,8'h00,8'h00,8'h00,8'h00,8'hd4,8'h24,8'h24,8'h24,8'h24,8'h91,8'hb6,8'h00,8'hfc,8'hfc,8'h6d,8'hb6,8'h91,8'h91,8'h91,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'h91,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00},
	{8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h36,8'h35,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'hfc,8'h6d,8'hda,8'hff,8'h00,8'h00,8'h6d,8'h24,8'h24,8'h6d,8'hb6,8'h91,8'h6d,8'hb6,8'hda,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'h91,8'h91,8'h90,8'hfc,8'h00,8'hb6,8'hb6,8'h91,8'h91,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8c,8'hd4,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hd4,8'h6d,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00},
	{8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h36,8'h7a,8'h7a,8'h7a,8'h7e,8'h7a,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'hfc,8'h00,8'hb6,8'hda,8'h00,8'h00,8'h6d,8'h00,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h6d,8'h6d,8'h00,8'h00,8'h00,8'h24,8'h24,8'h91,8'h91,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h00,8'hfc,8'hd4,8'hb6,8'h91,8'h91,8'h91,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd8,8'hfc,8'hf8,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00},
	{8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7e,8'h7a,8'h7e,8'h7e,8'h7e,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'hfc,8'h00,8'hb6,8'hb6,8'h00,8'h00,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h91,8'hfc,8'hfc,8'hb6,8'h00,8'h24,8'h24,8'hb6,8'hda,8'hda,8'hb6,8'hb6,8'hb6,8'hb6,8'h00,8'hfc,8'hfc,8'h6d,8'h91,8'h91,8'h91,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf8,8'hfc,8'hd4,8'hd4,8'hd4,8'hb0,8'hd8,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'hd4,8'hf8,8'hd4,8'hd4,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hda,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00},
	{8'h00,8'hff,8'hff,8'hff,8'hff,8'h36,8'h7a,8'h7a,8'h7e,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7a,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'hfc,8'h00,8'h6d,8'h91,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hfc,8'h36,8'h36,8'hdf,8'h36,8'hfc,8'h24,8'hb6,8'hb6,8'hff,8'hda,8'hda,8'hda,8'hb6,8'h00,8'hfc,8'hfc,8'h6d,8'h91,8'h91,8'h91,8'h91,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8c,8'hfc,8'hfc,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hd4,8'hd8,8'hd9,8'hb0,8'hb0,8'hb0,8'hb0,8'hd4,8'hf8,8'hf8,8'hd4,8'hf8,8'hf8,8'hd4,8'hf8,8'hf8,8'hd4,8'hd4,8'hd4,8'hb0,8'hda,8'hda,8'hda,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'hfc,8'h00,8'h6d,8'h91,8'h91,8'h91,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hfc,8'h36,8'h36,8'h9a,8'h36,8'h36,8'h35,8'hfd,8'hb6,8'h91,8'h91,8'hff,8'hda,8'hda,8'h00,8'hfc,8'hfc,8'h00,8'h91,8'h91,8'h91,8'h91,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb0,8'hfc,8'hfc,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hd9,8'hd8,8'hd4,8'hb0,8'hb0,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'hf8,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hda,8'hda,8'hda,8'hd4,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7e,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'hd8,8'h24,8'h00,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'h6d,8'hfc,8'h35,8'h36,8'hdf,8'h9a,8'h36,8'h9a,8'h9a,8'h9a,8'hfd,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h24,8'hfc,8'hfc,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hfc,8'hfc,8'hf8,8'hd8,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hf9,8'hd8,8'hd4,8'h90,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'hf8,8'hf8,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hda,8'hda,8'hda,8'hb0,8'hb0,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hff,8'hff,8'hff,8'hff,8'h36,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'hfc,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfc,8'h36,8'h36,8'hfd,8'h91,8'h00,8'h91,8'h91,8'h91,8'hfd,8'h9a,8'hb6,8'hb6,8'hb6,8'h91,8'h24,8'hfd,8'hfc,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hfc,8'hfc,8'hfc,8'hf8,8'hf9,8'hf9,8'hf8,8'hf8,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hfd,8'hf9,8'hfd,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hda,8'hda,8'hda,8'hb0,8'hb0,8'hb0,8'hb0,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7a,8'h7e,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h36,8'h36,8'h36,8'h36,8'h36,8'h35,8'h36,8'h36,8'h36,8'hfc,8'hd4,8'hf8,8'hfc,8'h36,8'h35,8'hb6,8'hb6,8'h00,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h9a,8'h9a,8'hd8,8'h00,8'hfc,8'hfd,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf8,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfe,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hfc,8'hd4,8'hd4,8'hd8,8'hd4,8'hd4,8'hd4,8'hd9,8'hfd,8'hfd,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hff,8'hda,8'hda,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7e,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'hfe,8'hb6,8'h91,8'h91,8'hff,8'hff,8'hff,8'hb6,8'h91,8'h91,8'hfd,8'h35,8'h35,8'h00,8'hfc,8'hd4,8'h24,8'h24,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hfc,8'hf8,8'hd4,8'hd4,8'hd8,8'hd4,8'hd4,8'hd4,8'hfd,8'hfd,8'hfc,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hda,8'hda,8'hda,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7e,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7a,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h35,8'hdf,8'hb6,8'hb6,8'hff,8'h91,8'h91,8'h91,8'h91,8'h91,8'hda,8'h6d,8'h00,8'h31,8'h00,8'hfc,8'hfc,8'h24,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hd4,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hfc,8'hfe,8'hfd,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hff,8'hff,8'hff,8'hb0,8'hb0,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7a,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'hdf,8'hfe,8'hb6,8'hff,8'hb6,8'hda,8'hb6,8'hb6,8'hb6,8'hb6,8'h24,8'h00,8'h00,8'hb0,8'hf8,8'hfc,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hff,8'hfe,8'hfc,8'hfc,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hd8,8'hd8,8'hd8,8'hd8,8'hd4,8'hf8,8'hfc,8'hfc,8'hfe,8'hfe,8'hfd,8'hfc,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'hf8,8'hd4,8'hd4,8'hd4,8'hff,8'hda,8'hd4,8'hb0,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h36,8'h36,8'h36,8'h36,8'h36,8'h35,8'hdf,8'hdf,8'hfe,8'hb6,8'hb6,8'hda,8'hb6,8'hda,8'h6d,8'h00,8'h00,8'h24,8'hfc,8'hf8,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfc,8'hfd,8'hfd,8'hfc,8'hfd,8'hfc,8'hfc,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfc,8'hfc,8'hf8,8'hd8,8'hf9,8'hd8,8'hf9,8'hd4,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hff,8'hff,8'hd4,8'hb0,8'hb0,8'hb0,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h76,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7a,8'h7e,8'h7a,8'h36,8'h36,8'h36,8'h36,8'hdf,8'hdf,8'hdf,8'hfe,8'hb6,8'hb6,8'hda,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hf8,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfc,8'hfc,8'hfd,8'hfc,8'hfc,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hf9,8'hf9,8'hf9,8'hd4,8'hfc,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfc,8'hf8,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'hf8,8'hd4,8'hd4,8'hd4,8'hda,8'hff,8'hff,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7a,8'h36,8'h36,8'h36,8'hdf,8'hdf,8'hdf,8'hdf,8'hfc,8'h24,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hfc,8'hf9,8'hd4,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'hd4,8'hff,8'hff,8'hda,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7e,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7a,8'h7e,8'h7e,8'h36,8'hff,8'hdf,8'hdf,8'hdf,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hd4,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfc,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hfc,8'hfd,8'hfc,8'hfd,8'hfd,8'hfc,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'hd4,8'hff,8'hff,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7a,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'hdf,8'hdf,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hb0,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hd9,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hf8,8'hf9,8'hf8,8'hf9,8'hf8,8'hf8,8'hd8,8'hf8,8'hf8,8'hd4,8'hff,8'hff,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hd4,8'hd4,8'hb0,8'hd9,8'hd9,8'hb6,8'hd9,8'hb6,8'hb6,8'hb6,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7e,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'hff,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfc,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hd9,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfe,8'hfe,8'hfe,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hd8,8'hd4,8'hff,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hd4,8'hb0,8'hda,8'hda,8'hda,8'hda,8'hd9,8'hd4,8'hd9,8'hb6,8'hb6,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7b,8'h7e,8'h7e,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hb0,8'hfc,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hff,8'hfe,8'hfe,8'hff,8'hfd,8'hfe,8'hfd,8'hfd,8'hfe,8'hfd,8'hfe,8'hfe,8'hfd,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hd9,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hff,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hfd,8'hfc,8'hf8,8'hf9,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'hff,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hda,8'hda,8'hd9,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hda,8'hff,8'hff,8'h7a,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hd4,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfd,8'hfc,8'hfc,8'hfc,8'hfd,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfc,8'hfd,8'hf9,8'hfc,8'hf9,8'hf8,8'hd8,8'hd8,8'hf8,8'hff,8'hd8,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hda,8'hda,8'hda,8'hd4,8'hb0,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb0,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hda,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7b,8'h7b,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfc,8'hfc,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hb6,8'hb6,8'hda,8'hda,8'hff,8'hff,8'hda,8'hfe,8'hfd,8'hfd,8'hfd,8'hfc,8'hf9,8'hf9,8'hf9,8'hf8,8'hf9,8'hf9,8'hff,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hda,8'hda,8'hd4,8'hd4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7a,8'h7e,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7b,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h00,8'h00,8'h24,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hb0,8'hfc,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfd,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hb6,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'hb6,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hf9,8'hf9,8'hf9,8'hf8,8'hf8,8'hd8,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hfd,8'hfd,8'hda,8'hd4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hda,8'hda,8'hff,8'hff,8'h76,8'h7a,8'h7b,8'h7b,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hb0,8'hfc,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hb6,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hf9,8'hf9,8'hf8,8'hf8,8'hd8,8'hf8,8'hd8,8'hd8,8'hd4,8'hd8,8'hd4,8'hd4,8'hd4,8'hda,8'hda,8'hd4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hff,8'hff,8'hff,8'hff,8'hff,8'h7a,8'h7a,8'h7e,8'h7b,8'h7e,8'h7e,8'h7e,8'h7e,8'h36,8'h36,8'h7e,8'h7e,8'h7e,8'h7b,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hfc,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hff,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hda,8'hff,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'h91,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hf9,8'hf8,8'hf9,8'hf8,8'hd8,8'hd4,8'hd4,8'hd8,8'hd8,8'hd4,8'hfd,8'hda,8'hd4,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hff,8'hda,8'hda,8'hff,8'h7a,8'h7a,8'h76,8'h7b,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h00,8'h00,8'h8c,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hff,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hb6,8'hfd,8'hfd,8'hfd,8'hfd,8'hf8,8'hf9,8'hf9,8'hf9,8'hf9,8'hd8,8'hd8,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hda,8'hda,8'hd4,8'h00,8'h24,8'h91,8'h91,8'h91,8'h91,8'h91,8'h00,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h7a,8'h7a,8'h7a,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7e,8'h7b,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hb0,8'hfc,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hff,8'hfe,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hd9,8'hfd,8'hfd,8'hfd,8'hfc,8'hfd,8'hf9,8'hf9,8'hf9,8'hf9,8'hd8,8'hf8,8'hd4,8'hd4,8'hd4,8'hda,8'hda,8'hd9,8'h6d,8'hb6,8'h91,8'h91,8'hb6,8'h91,8'h91,8'h91,8'h91,8'h91,8'h6d,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h7a,8'h7a,8'h76,8'h7e,8'h7e,8'h7e,8'h7b,8'h7e,8'h7e,8'h7e,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hb0,8'hfc,8'hfc,8'hff,8'hfe,8'hff,8'hfe,8'hff,8'hfe,8'hfe,8'hff,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdf,8'hda,8'hda,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hf8,8'hf9,8'hf8,8'hd4,8'hd4,8'hd4,8'hda,8'hda,8'hd4,8'h91,8'h6d,8'h00,8'h00,8'h00,8'hb6,8'h91,8'h91,8'h91,8'h91,8'h6d,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h32,8'h35,8'h36,8'h7a,8'h7e,8'h7b,8'h7e,8'h7e,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hb0,8'hfc,8'hfc,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hb6,8'hd9,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hf9,8'hf9,8'hf9,8'hf9,8'hf9,8'hd8,8'hd8,8'hd8,8'hd8,8'hfd,8'hfd,8'hd4,8'h00,8'h00,8'h91,8'h00,8'h00,8'h00,8'h00,8'h91,8'h91,8'h91,8'h91,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h35,8'h35,8'h32,8'h36,8'h36,8'h7b,8'h7e,8'h00,8'h00,8'h24,8'h24,8'h6d,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hb0,8'hfc,8'hfc,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hb6,8'hda,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hf9,8'hf9,8'hd8,8'hd8,8'hd8,8'hd8,8'hd4,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h91,8'h91,8'h91,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h35,8'h32,8'h35,8'h35,8'h36,8'h36,8'h00,8'h00,8'h24,8'h24,8'hff,8'h24,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hb0,8'hfc,8'hfc,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hb6,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hf9,8'hf8,8'hd8,8'hd8,8'hd4,8'hd9,8'hfd,8'hd4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h91,8'h91,8'h91,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h35,8'h35,8'h36,8'h35,8'h36,8'h00,8'h00,8'h24,8'h24,8'hff,8'hff,8'h24,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hfd,8'hf9,8'hf9,8'hf8,8'hd8,8'hd8,8'hda,8'hda,8'hd8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h91,8'h91,8'h91,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h35,8'h32,8'h35,8'h35,8'h00,8'h00,8'h24,8'h24,8'hff,8'hff,8'hff,8'h24,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hfd,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfd,8'hf9,8'hf9,8'hf8,8'hd8,8'hd8,8'hd4,8'hda,8'hda,8'hd8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h91,8'h91,8'hb6,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h35,8'h35,8'h32,8'h36,8'h00,8'h24,8'h24,8'hff,8'hff,8'hff,8'h24,8'hd4,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hfd,8'hfe,8'hfd,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hfd,8'hf9,8'hf9,8'hf8,8'hf8,8'hd8,8'hda,8'hda,8'hd4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h91,8'hda,8'h91,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h35,8'h36,8'h36,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'h24,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hb6,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hfd,8'hfd,8'hf9,8'hf8,8'hd8,8'hd8,8'hda,8'hd8,8'hd9,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hda,8'hda,8'h91,8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h7a,8'h76,8'h7e,8'h00,8'h24,8'hb6,8'hff,8'hff,8'hff,8'hff,8'h24,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hf9,8'hd8,8'hd8,8'hfd,8'hd4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hda,8'hda,8'h91,8'h24,8'hff,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h7a,8'h76,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'h91,8'h24,8'hfc,8'hfc,8'hf8,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hf9,8'hf9,8'hf9,8'hd8,8'hda,8'hd4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hda,8'hda,8'hda,8'h00,8'h24,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h7a,8'h7a,8'h00,8'h24,8'h6d,8'hff,8'hff,8'hff,8'hff,8'h24,8'hfc,8'hfc,8'hb0,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hf9,8'hd8,8'hd8,8'hfd,8'hd8,8'h00,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hb6,8'hb6,8'hda,8'hda,8'h6d,8'h00,8'h24,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h76,8'h7a,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'h24,8'h24,8'hfc,8'hb0,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hf9,8'hd8,8'hd8,8'hda,8'hd8,8'h00,8'hb6,8'hb6,8'h00,8'h00,8'h91,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h24,8'h24,8'h24,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h7a,8'h00,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'h24,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hda,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hd4,8'hf9,8'hf9,8'hd8,8'hd8,8'hda,8'hd8,8'h00,8'hb6,8'hb6,8'hb6,8'h24,8'hb6,8'hb6,8'hb6,8'h00,8'h91,8'h91,8'h24,8'h24,8'h24,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h7a,8'h00,8'h24,8'hb6,8'hff,8'hff,8'hff,8'h24,8'h24,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfd,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hd9,8'hf9,8'hf9,8'hd8,8'hd8,8'hd8,8'hd8,8'hda,8'hd4,8'h24,8'hb6,8'hb6,8'hff,8'hff,8'hb6,8'hda,8'h00,8'h00,8'h91,8'h91,8'h24,8'hda,8'h00,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h76,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'h24,8'hfc,8'hb0,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hd8,8'hd8,8'hd8,8'hd4,8'hda,8'hd4,8'h00,8'h24,8'hff,8'hff,8'hff,8'hff,8'h24,8'h00,8'h24,8'h91,8'h91,8'hda,8'hda,8'h00,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff},
	{8'hda,8'hda,8'hdf,8'hda,8'hff,8'h7a,8'h00,8'h24,8'hff,8'hff,8'hff,8'h24,8'h24,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hd9,8'hd8,8'hd8,8'hd8,8'hd8,8'hda,8'hd8,8'h00,8'h6d,8'hda,8'hff,8'hff,8'h91,8'h00,8'h00,8'h91,8'h91,8'hda,8'hda,8'hda,8'h24,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h00,8'h00,8'h24,8'hff,8'hff,8'h91,8'h24,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hda,8'hfe,8'hfe,8'hfd,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hd9,8'hf9,8'hf9,8'hf9,8'hf9,8'hd8,8'hd8,8'hda,8'hd8,8'h91,8'hda,8'hda,8'hda,8'h91,8'h91,8'h91,8'h00,8'h91,8'hff,8'hda,8'h24,8'h24,8'h24,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h00,8'hd4,8'h24,8'hff,8'hff,8'h24,8'hfc,8'hb0,8'hfc,8'hfc,8'hfc,8'hfc,8'hfe,8'hfd,8'hfd,8'hfd,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hd9,8'hf9,8'hd9,8'hf9,8'hd8,8'hd8,8'hda,8'hff,8'hda,8'hda,8'hda,8'h24,8'h24,8'h91,8'h91,8'h91,8'hda,8'hda,8'h6d,8'h00,8'h00,8'h24,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h00,8'hfc,8'h24,8'hff,8'h24,8'h24,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hd9,8'hf9,8'hf9,8'hd8,8'hd9,8'hd8,8'hd8,8'hff,8'hfe,8'hda,8'hda,8'h00,8'h24,8'h24,8'h24,8'h91,8'hda,8'hda,8'h24,8'h24,8'h6d,8'h6d,8'h24,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'h00,8'h00,8'hfc,8'h24,8'h6d,8'h24,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hff,8'hfe,8'hff,8'hfe,8'hff,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hd8,8'hd8,8'hd8,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'h00,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h24,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'h00,8'hfc,8'hfc,8'h24,8'h24,8'hfc,8'hf8,8'hfc,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hd9,8'hf9,8'hd8,8'hd9,8'hd8,8'hff,8'hff,8'hff,8'hfe,8'hd4,8'h00,8'h00,8'h00,8'h00,8'hda,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h24,8'hda,8'hb6,8'hb6,8'hb6,8'hda,8'hda,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'h00,8'hfc,8'hfc,8'hfc,8'h24,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hb0,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hd4,8'hd4,8'hd8,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hda,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hd8,8'hd8,8'hff,8'hff,8'hff,8'hd8,8'hd4,8'hd4,8'h00,8'h00,8'h00,8'hff,8'h00,8'h00,8'h91,8'h24,8'h00,8'h24,8'h24,8'h00,8'h24,8'hda,8'hda,8'hda,8'hb6,8'hb6,8'hda,8'hff},
	{8'hb6,8'hda,8'hda,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'h6d,8'h90,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hd4,8'hb0,8'hb0,8'h90,8'hb0,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hd4,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hd8,8'hd8,8'hff,8'hff,8'hff,8'hd8,8'hd8,8'hd4,8'hb0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h91,8'h91,8'h00,8'h00,8'h6d,8'h00,8'h24,8'hda,8'hda,8'hb6,8'hb6,8'hb6,8'hda,8'hff},
	{8'hda,8'hda,8'hda,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'h00,8'h6d,8'h24,8'h24,8'h90,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hb0,8'hb0,8'h6d,8'h6d,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hda,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hfe,8'hfe,8'hfd,8'hd9,8'hfd,8'hf9,8'hfd,8'hf9,8'hd8,8'hff,8'hff,8'hff,8'hd4,8'hd4,8'hd8,8'hb0,8'hb0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h6d,8'h91,8'h24,8'h6d,8'h6d,8'h00,8'h24,8'hda,8'hb6,8'hb6,8'hb6,8'hb6,8'hda,8'hff},
	{8'hda,8'hb6,8'h91,8'h00,8'hfc,8'hfc,8'hfc,8'hf8,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h90,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hb0,8'hb0,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hda,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hff,8'hff,8'hff,8'hd4,8'hd4,8'hd4,8'hb0,8'hd9,8'hb0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h91,8'h00,8'h00,8'h24,8'h6d,8'h00,8'h24,8'hb6,8'hda,8'hda,8'hda,8'hb6,8'hda,8'hff},
	{8'hb6,8'hda,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'h8c,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h8c,8'hb0,8'hb0,8'h90,8'h90,8'hb0,8'hb0,8'h90,8'h8c,8'h90,8'h90,8'h8c,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h00,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'hd4,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfd,8'hda,8'hfe,8'hfe,8'hfe,8'hfe,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfe,8'hfd,8'hfd,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hf9,8'hf9,8'hff,8'hff,8'hff,8'hd4,8'hd8,8'hd4,8'hd4,8'hd4,8'hda,8'hb0,8'h00,8'h00,8'h00,8'h00,8'h91,8'h91,8'h91,8'h00,8'h00,8'h24,8'h6d,8'h6d,8'h24,8'hda,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'hda,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hda,8'hfd,8'hfd,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfd,8'hfd,8'hfd,8'hd9,8'hff,8'hff,8'hff,8'hd8,8'hd8,8'hd8,8'hd4,8'hb0,8'hb0,8'hd4,8'hb0,8'h00,8'h00,8'h00,8'h00,8'h91,8'h91,8'h00,8'h00,8'h00,8'h24,8'h6d,8'h6d,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'hb6,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hff,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hd9,8'hff,8'hff,8'hff,8'hfd,8'hd8,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'h90,8'h00,8'h00,8'h24,8'h6d,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hb6,8'hda,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h00,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'hf9,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hff,8'hff,8'hff,8'hfd,8'hd8,8'hd8,8'hd4,8'hd4,8'hd9,8'hb0,8'hd4,8'hb0,8'hb0,8'h90,8'hb0,8'h00,8'h24,8'h91,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h6d,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hff,8'h00,8'h8c,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h00,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hff,8'hff,8'hff,8'hfd,8'hf9,8'hd8,8'hd4,8'hd9,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'h90,8'h91,8'h91,8'h91,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'h00,8'hfc,8'hfc,8'hfc,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h8c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h00,8'hb0,8'hfc,8'hfc,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hff,8'hff,8'hff,8'hf9,8'hd9,8'hd9,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hd4,8'hb0,8'hb0,8'h90,8'h90,8'h00,8'h91,8'h6d,8'h24,8'h24,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'h00,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h90,8'h90,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h90,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hff,8'hff,8'hfd,8'hf9,8'hd8,8'hd8,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'h90,8'h90,8'h00,8'h91,8'h91,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'h00,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hd4,8'h90,8'h90,8'h8c,8'h8c,8'h90,8'h90,8'h8c,8'h90,8'hd4,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'h91,8'h91,8'hb6,8'hb6,8'hb6,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hff,8'hff,8'hd8,8'hd8,8'hd8,8'hd8,8'hd8,8'hd4,8'hd9,8'hd4,8'hd4,8'hb0,8'hb0,8'hd4,8'hb0,8'hb0,8'h90,8'h90,8'h90,8'h8c,8'h91,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'h00,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfc,8'hfd,8'hfc,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hb6,8'h91,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h91,8'h91,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hff,8'hff,8'hf9,8'hd8,8'hf9,8'hd8,8'hd8,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'h90,8'h90,8'h90,8'h90,8'h90,8'h91,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'h00,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfc,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'hfd,8'hfd,8'hfe,8'h91,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'hb6,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h6d,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hff,8'hff,8'hf9,8'hf9,8'hd8,8'hd8,8'hd8,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd9,8'h91,8'hd4,8'hb0,8'hb0,8'hb0,8'h90,8'h90,8'h90,8'h90,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'h00,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hfd,8'hfc,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'hfe,8'hfe,8'hfd,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'hfd,8'hfd,8'hfd,8'hf9,8'hff,8'hff,8'hf9,8'hd8,8'hd8,8'hd8,8'hd8,8'hd4,8'hd4,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hd4,8'h90,8'hb0,8'h90,8'h90,8'h90,8'h8c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'h00,8'h00,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hfd,8'hfd,8'hfc,8'hfd,8'hfc,8'hfc,8'hfc,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfc,8'hfd,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfe,8'hfe,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'h6d,8'h91,8'h91,8'h91,8'h6d,8'h91,8'h91,8'hb6,8'hb6,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hfd,8'hf9,8'hff,8'hff,8'hf9,8'hf9,8'hf9,8'hd8,8'hd9,8'hd9,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'h90,8'h90,8'h90,8'h90,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'hda,8'h00,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'h24,8'h91,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'h91,8'h6d,8'h91,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h6d,8'h6d,8'h6d,8'h24,8'hff,8'hff,8'hfd,8'hd8,8'hf9,8'hd8,8'hd8,8'hd8,8'hd8,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hd4,8'hb0,8'hb0,8'h90,8'h90,8'h90,8'h90,8'h90,8'h8c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'hda,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfc,8'hfd,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf9,8'h00,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h91,8'h91,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h6d,8'h24,8'h6d,8'hff,8'hff,8'hd8,8'hf9,8'hd8,8'hd8,8'hd8,8'hd8,8'hd8,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h91,8'h90,8'h90,8'h90,8'h90,8'h8c,8'h90,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'hda,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfc,8'hfd,8'hfc,8'hfc,8'hfc,8'hfd,8'hfc,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h91,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h91,8'h6d,8'h24,8'hff,8'hff,8'hf8,8'hd8,8'hf9,8'hd8,8'hd8,8'hd4,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'h90,8'h90,8'h90,8'h90,8'h8c,8'h8c,8'h90,8'h6d,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'hda,8'h00,8'h00,8'hfc,8'hd4,8'hd4,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfd,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h91,8'h6d,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'hff,8'h6d,8'h24,8'hf9,8'hf8,8'hd8,8'hd8,8'hd8,8'hd8,8'hd4,8'hd8,8'hd4,8'hd8,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'h90,8'h90,8'h8c,8'h8c,8'h8c,8'h8c,8'h00,8'h00,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'hda,8'h6d,8'h00,8'hfc,8'hfc,8'hd4,8'hd4,8'hd4,8'hd4,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfd,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h24,8'h24,8'h24,8'hd8,8'hd8,8'hd8,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'h90,8'h90,8'h8c,8'h90,8'h90,8'h8c,8'h8c,8'h8c,8'h8c,8'h00,8'h00,8'h00,8'h6d,8'h24,8'h24,8'h6d,8'h24,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'hda,8'hda,8'h00,8'hfc,8'hfc,8'hfc,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h91,8'h91,8'h91,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h6d,8'h24,8'h24,8'h24,8'hd8,8'hd8,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd8,8'hd4,8'hd4,8'hb0,8'hb0,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'h8c,8'h90,8'h90,8'h8c,8'h8c,8'h90,8'h8c,8'h8c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hda,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'hda,8'hda,8'h00,8'hfc,8'hfc,8'hfc,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hd4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h91,8'h91,8'h6d,8'h91,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h6d,8'h24,8'h00,8'h24,8'hd4,8'hd8,8'hd4,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'h24,8'h90,8'h90,8'h90,8'h8c,8'h8c,8'h8c,8'h8c,8'h8c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'hda,8'hda,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h6d,8'h91,8'h91,8'h91,8'h6d,8'h91,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h24,8'h6d,8'h24,8'h6d,8'h91,8'h91,8'h91,8'h91,8'h91,8'h24,8'h24,8'h00,8'h00,8'h00,8'hd8,8'hd4,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h8c,8'h90,8'h90,8'h90,8'h90,8'h8c,8'h90,8'h8c,8'h8c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'h00,8'hfc,8'hfc,8'hfc,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd8,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'hd4,8'hd4,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h24,8'h24,8'hff,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'hd8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'h24,8'hb0,8'h90,8'h90,8'h90,8'h90,8'h8c,8'h90,8'h8c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h2d,8'h2d,8'h24,8'h24,8'hda,8'hda,8'hb6,8'hb6,8'hb6,8'hda,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'h00,8'hf8,8'hfc,8'hfc,8'hfc,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h00,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'h8c,8'h90,8'h90,8'h90,8'h90,8'h90,8'h8c,8'h8c,8'h8c,8'h90,8'h00,8'h00,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h31,8'h00,8'h24,8'hda,8'hda,8'hb6,8'hb6,8'hb6,8'hda,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h00,8'h24,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'h24,8'hb0,8'hb0,8'h90,8'h90,8'h90,8'h8c,8'h90,8'h8c,8'h8c,8'h00,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h31,8'h2d,8'h2d,8'h2d,8'h24,8'hda,8'hb6,8'hda,8'hb6,8'hb6,8'hb6,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hd4,8'hfc,8'h24,8'h24,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hd4,8'hb0,8'hb0,8'h8c,8'h90,8'h90,8'h90,8'h90,8'h90,8'h8c,8'h90,8'h90,8'h8c,8'h00,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h31,8'h00,8'h24,8'hda,8'hb6,8'hda,8'hda,8'hb6,8'hda,8'hff},
	{8'hda,8'hda,8'hda,8'hda,8'hff,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hd4,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'h8c,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hd4,8'hb0,8'hb0,8'hb0,8'h8c,8'hb0,8'hb0,8'h90,8'hb0,8'h90,8'h90,8'h8c,8'h90,8'h8c,8'h90,8'h00,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h31,8'h2d,8'h2d,8'h2d,8'h00,8'h24,8'hb6,8'hb6,8'hb6,8'hb6,8'hda,8'hb6,8'hff},
	{8'hff,8'hda,8'hda,8'hda,8'hff,8'h7b,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hd4,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hd4,8'hb0,8'hb0,8'hb0,8'h8c,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'h90,8'h90,8'h8c,8'h8c,8'h8c,8'h00,8'h2d,8'h2d,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h2d,8'h24,8'hb6,8'hb6,8'hb6,8'hda,8'hb6,8'hb6,8'hff},
	{8'hff,8'hda,8'hda,8'hda,8'hff,8'h76,8'h7b,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb0,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hd4,8'hb0,8'h8c,8'hb0,8'hb0,8'hb0,8'h90,8'hb0,8'hb0,8'h90,8'h90,8'h90,8'h8c,8'h8c,8'h00,8'h2d,8'h2d,8'h2d,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h31,8'h32,8'h76,8'h2d,8'h24,8'hb6,8'hda,8'hb6,8'hda,8'hda,8'hb6,8'h00},
	{8'h00,8'hda,8'hda,8'hda,8'hff,8'hdf,8'h7b,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h24,8'hfc,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'hd4,8'hd4,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8c,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'h8c,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'hb0,8'hb0,8'hb0,8'h90,8'h8c,8'h90,8'h90,8'h00,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h76,8'h76,8'h76,8'h76,8'h2d,8'h24,8'hb6,8'hda,8'hda,8'hb6,8'hda,8'hb6,8'h00},
	{8'h00,8'hda,8'hda,8'hda,8'hff,8'hff,8'h7b,8'h7b,8'h00,8'h24,8'hfc,8'hfc,8'hfc,8'hfc,8'hd4,8'hfc,8'hfc,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfc,8'hd4,8'hb0,8'hd4,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'h8c,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'h90,8'h90,8'h8c,8'h90,8'h00,8'h2d,8'h24,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h31,8'h2d,8'h2d,8'h7b,8'h76,8'h76,8'h32,8'h76,8'h2d,8'h24,8'hb6,8'hb6,8'hda,8'hda,8'hb6,8'hb6,8'h00},
	{8'h00,8'hda,8'hda,8'hda,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h00,8'h90,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb0,8'hd4,8'hd4,8'hd4,8'h8c,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'h90,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'hb0,8'h90,8'h90,8'h90,8'h00,8'h00,8'h31,8'h31,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h31,8'h31,8'h31,8'h7b,8'h7b,8'h7b,8'h76,8'h76,8'h32,8'h2d,8'h24,8'hda,8'hda,8'hda,8'hda,8'hb6,8'hda,8'h00},
	{8'h00,8'hda,8'hda,8'hda,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'hd4,8'hd4,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'hb0,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hd4,8'hd4,8'hb0,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'hb0,8'hb0,8'h90,8'h90,8'h00,8'h00,8'h2d,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h2d,8'h31,8'h31,8'h31,8'h7b,8'h7b,8'h7b,8'h7b,8'h76,8'h76,8'h32,8'h2d,8'h24,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00},
	{8'h00,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h31,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hd4,8'hd4,8'hd4,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'hb0,8'hf8,8'hd4,8'hd4,8'hd4,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'h90,8'h00,8'h31,8'h2d,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h7b,8'h7b,8'h76,8'h7b,8'h7b,8'h76,8'h76,8'h32,8'h2d,8'h24,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00},
	{8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h31,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hb0,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'hfc,8'hd4,8'hd4,8'hd4,8'hd4,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h8c,8'hfc,8'hf8,8'hfc,8'hf8,8'hf8,8'hf8,8'hd4,8'hd4,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h00,8'h00,8'h31,8'h31,8'h31,8'h24,8'h2d,8'h31,8'h31,8'h31,8'h2d,8'h31,8'h2d,8'h7b,8'h7b,8'h7b,8'h76,8'h7b,8'h76,8'h76,8'h76,8'h32,8'h2d,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00},
	{8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h31,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'hf8,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb0,8'h90,8'h24,8'h00,8'h00,8'h31,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h7b,8'h7b,8'h7b,8'h7b,8'h76,8'h7b,8'h76,8'h76,8'h32,8'h31,8'h24,8'hb6,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00},
	{8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h31,8'h31,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'hb0,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'hf8,8'hfc,8'hf8,8'hfc,8'hf8,8'hfc,8'hfc,8'hf8,8'hf8,8'hd4,8'hf8,8'hd4,8'hf8,8'hd4,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'hb0,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'h00,8'h00,8'h31,8'h31,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h31,8'h31,8'h31,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h76,8'h76,8'h76,8'h76,8'h2d,8'h24,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00},
	{8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h31,8'h32,8'h32,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hd4,8'hd4,8'hb0,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'hfc,8'hf8,8'hfc,8'hf8,8'hfc,8'hf8,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hd4,8'hd4,8'hb0,8'hd4,8'hd4,8'hb0,8'hb0,8'h00,8'h00,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h76,8'h76,8'h76,8'h76,8'h32,8'h2d,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h31,8'h31,8'h32,8'h32,8'h00,8'h00,8'h00,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hfc,8'hfc,8'hf8,8'hf8,8'hf8,8'hfc,8'hfc,8'hf8,8'hf8,8'hf8,8'hf8,8'hd4,8'h00,8'h00,8'hd4,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hb0,8'hb0,8'h00,8'h00,8'h00,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h32,8'h76,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h76,8'h76,8'h76,8'h76,8'h2d,8'h24,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h31,8'h31,8'h31,8'h31,8'h32,8'h00,8'h00,8'h00,8'h00,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hf8,8'hfc,8'hfc,8'h8c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd4,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hb0,8'hd4,8'hd4,8'h00,8'h00,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h7b,8'h76,8'h32,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h76,8'h76,8'h76,8'h32,8'h2d,8'hb6,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h31,8'h32,8'h31,8'h32,8'h2d,8'h2d,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'hfc,8'hfc,8'hfc,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h00,8'hf8,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'hd4,8'h90,8'h00,8'h00,8'h00,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h7b,8'h7b,8'h7b,8'h7b,8'h32,8'h76,8'h7b,8'h7b,8'h7b,8'h76,8'h76,8'h76,8'h76,8'h76,8'h2d,8'h91,8'hda,8'hda,8'hda,8'hda,8'hdf,8'hda,8'hff,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h32,8'h32,8'h31,8'h2d,8'h2d,8'h2d,8'h2d,8'h31,8'h31,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h90,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hfc,8'hf8,8'h8c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h32,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h00,8'h8c,8'hf8,8'hf8,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h32,8'h7b,8'h7b,8'h76,8'h7b,8'h7b,8'h76,8'h76,8'h2d,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h31,8'h2d,8'h2d,8'h2d,8'h31,8'h32,8'h31,8'h2d,8'h2d,8'h2d,8'h2d,8'h31,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h31,8'h32,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h76,8'h76,8'h76,8'h76,8'h2d,8'h91,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h32,8'h31,8'h31,8'h32,8'h31,8'h2d,8'h2d,8'h2d,8'h31,8'h32,8'h32,8'h31,8'h32,8'h31,8'h31,8'h31,8'h31,8'h31,8'h32,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h32,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h76,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h76,8'h76,8'h76,8'h2d,8'hb6,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h2d,8'h31,8'h32,8'h31,8'h32,8'h31,8'h31,8'h31,8'h31,8'h31,8'h32,8'h31,8'h32,8'h32,8'h31,8'h32,8'h31,8'h31,8'h31,8'h32,8'h31,8'h31,8'h31,8'h31,8'h31,8'h32,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h24,8'h31,8'h31,8'h31,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h76,8'h7b,8'h7b,8'h76,8'h76,8'h76,8'h76,8'h91,8'hda,8'hff,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h2d,8'h2d,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h31,8'h32,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h32,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h31,8'h76,8'h76,8'h76,8'h7b,8'h31,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h76,8'h7b,8'h76,8'h76,8'h7b,8'h7b,8'h7b,8'h76,8'h76,8'h7b,8'h76,8'h76,8'h76,8'h32,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h32,8'h76,8'h7b,8'h31,8'h32,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h32,8'h31,8'h31,8'h31,8'h31,8'h32,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h76,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h32,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h76,8'h7b,8'h76,8'h76,8'h7b,8'h7b,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h32,8'h76,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h76,8'h2d,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h31,8'h2d,8'h32,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h76,8'h31,8'h31,8'h2d,8'h31,8'h31,8'h31,8'h7b,8'h7b,8'h76,8'h7b,8'h76,8'h76,8'h7b,8'h76,8'h7b,8'h76,8'h7b,8'h7b,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h32,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdf,8'h7b,8'h7b,8'h76,8'h32,8'h32,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h7b,8'h76,8'h7b,8'h7b,8'h7b,8'h7b,8'h76,8'h76,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h32,8'h76,8'h7b,8'h7b,8'h7b,8'h76,8'h76,8'h7b,8'h76,8'h76,8'h76,8'h76,8'h76,8'h7b,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h76,8'h32,8'h76,8'h76,8'h76,8'h76,8'h76,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'hff,8'hda,8'hda,8'hda,8'hda,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hda,8'hff,8'hff,8'hff,8'hff,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'hff,8'hda,8'hda,8'hda,8'hda,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hda,8'hda,8'hda,8'hda,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hda,8'hda,8'hff,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hff,8'hda,8'hff,8'hff,8'hff,8'hda,8'hff,8'hff,8'hff,8'hda,8'hff,8'hff,8'hda,8'hda,8'hff,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hff,8'hda,8'hff,8'hda,8'hff,8'hda,8'hda,8'hff,8'hda,8'hff,8'hda,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hff,8'hda,8'hff,8'hda,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'hff,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'hda,8'hff,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hda,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}};

 
 
//////////--------------------------------------------------------------------------------------------------------------= 
always_ff@(posedge clk or negedge resetN) 
begin 
	if(!resetN)  
		RGBout <= object_colors[offsetY][offsetX]; 	
	else begin 
		RGBout <= TRANSPARENT_ENCODING ; // default   
		if (InsideRectangle == 1'b1) 
			RGBout <= object_colors[offsetY][offsetX]; 		 
	end 
end 
 
//////////--------------------------------------------------------------------------------------------------------------= 
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
 
endmodule 
