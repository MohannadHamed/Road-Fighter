
 module gameOverBitMap (

					input	logic	clk, 
					input	logic	resetN, 
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY, 
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input	logic	gameOver, //input that the pixel is within a bracket 
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ; 
 
 
// generating the bitmap 
 

localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel  
logic[0:63][0:63][7:0] object_colors = {
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hcd,8'ha4,8'had,8'hcd,8'hc5,8'ha4,8'ha5,8'hcd,8'ha4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha4,8'ha4,8'had,8'hc4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha4,8'ha4,8'ha4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha4,8'hc4,8'hc5,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha4,8'ha4,8'hcd,8'hc5,8'hcd,8'hc5,8'ha5,8'ha4,8'ha4,8'hcd,8'h60,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'he4,8'hf1,8'hf1,8'hf1,8'hf1,8'hf1,8'hf2,8'hf1,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'he0,8'hec,8'he4,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'he4,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'he0,8'hed,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h00,8'he0,8'hf1,8'hf1,8'hf1,8'hf1,8'hf1,8'hf1,8'hf1,8'hf1,8'he4,8'h60,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'he0,8'hed,8'he4,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'hc0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'he0,8'he4,8'he4,8'h80,8'h80,8'he4,8'he4,8'hed,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'he4,8'hf1,8'hc0,8'h00,8'h00,8'h00,8'hec,8'he4,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'h60,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h80,8'hc0,8'h80,8'h60,8'h60,8'h60,8'h60,8'h60,8'h60,8'h60,8'h60,8'h00,8'h00,8'h00,8'h00,8'h00,8'h60,8'he4,8'he0,8'h80,8'h20,8'h60,8'ha0,8'he0,8'he4,8'h60,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'he0,8'he0,8'he4,8'h60,8'h60,8'h60,8'he0,8'he0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'he0,8'h80,8'h60,8'h60,8'h60,8'h60,8'h60,8'h60,8'h20,8'h20,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h80,8'ha0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'he0,8'he4,8'h80,8'h80,8'h00,8'h00,8'h80,8'h80,8'he4,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h80,8'ha0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'hc0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h80,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h80,8'h80,8'he0,8'he0,8'h80,8'h80,8'h80,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h80,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h80,8'he0,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'h80,8'h80,8'h80,8'h80,8'hc0,8'h80,8'h80,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h80,8'hc0,8'hc0,8'h00,8'h00,8'he0,8'hed,8'he4,8'he4,8'he4,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'hc0,8'h00,8'h00,8'h00,8'h00,8'hc0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'he0,8'h80,8'h00,8'h00,8'ha0,8'ha0,8'h80,8'h00,8'h80,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'hec,8'he4,8'hed,8'hed,8'hed,8'hed,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h80,8'hc0,8'ha0,8'h00,8'h00,8'hc0,8'h80,8'he0,8'ha0,8'he0,8'he4,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'h80,8'h00,8'h00,8'h80,8'ha0,8'h80,8'h00,8'h80,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'he0,8'ha0,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h80,8'hc0,8'hc0,8'h00,8'h00,8'h80,8'h80,8'h80,8'h80,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'h80,8'h00,8'h00,8'h80,8'h80,8'h80,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'he0,8'h80,8'h60,8'h80,8'h80,8'h80,8'h80,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h80,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'h80,8'h80,8'h80,8'h80,8'ha0,8'h80,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'ha0,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h80,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h80,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h80,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'ha0,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h80,8'ha0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'h80,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'he4,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'he0,8'he0,8'he0,8'hec,8'he0,8'he4,8'he0,8'he4,8'ha4,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h80,8'h80,8'ha0,8'he0,8'he0,8'he0,8'he4,8'he0,8'he0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'h80,8'h00,8'h00,8'h00,8'h00,8'hc0,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'h60,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'he4,8'h80,8'h80,8'h80,8'h80,8'ha0,8'h80,8'h80,8'he4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'h80,8'h80,8'h00,8'h00,8'h00,8'h00,8'h80,8'ha0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'h80,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'h80,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'h80,8'ha0,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'h60,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'he0,8'he0,8'h20,8'h00,8'h00,8'h00,8'h00,8'he0,8'he0,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'he0,8'he0,8'he4,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'h00,8'h00,8'h00,8'h00,8'h80,8'ha0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'ha0,8'he0,8'h80,8'h80,8'h80,8'hc0,8'h80,8'h80,8'he4,8'he0,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h80,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'he0,8'hc0,8'ha0,8'ha0,8'h80,8'h80,8'h80,8'ha0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h80,8'h80,8'ha0,8'h80,8'h80,8'hc0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h80,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h80,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h80,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h80,8'hc0,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'h80,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h80,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'he0,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'hc0,8'h80,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h80,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h80,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'h80,8'h80,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h80,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he4,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'h80,8'h80,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h80,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'hc0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h80,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'he4,8'he0,8'hc4,8'ha0,8'hc0,8'hc0,8'hc0,8'he4,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'he0,8'he0,8'hec,8'he0,8'he0,8'he0,8'he0,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'ha0,8'hc0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h80,8'hc0,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'hc0,8'h80,8'h80,8'h80,8'h80,8'ha0,8'he0,8'he0,8'he0,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h80,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h80,8'ha0,8'he0,8'h20,8'h00,8'h00,8'h00,8'h00,8'he0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h80,8'h80,8'he0,8'h80,8'h80,8'h80,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h80,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h80,8'h80,8'h80,8'he0,8'he0,8'h00,8'h00,8'he0,8'he0,8'h80,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'he0,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'h80,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h80,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'h80,8'he0,8'he0,8'he0,8'he0,8'ha0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'ha0,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h80,8'he0,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'he0,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'h80,8'ha0,8'he0,8'he0,8'ha0,8'h80,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'h80,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h80,8'h80,8'hc0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hc0,8'h80,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h60,8'h80,8'h80,8'h80,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'he0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'hc0,8'h80,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'ha0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'ha0,8'ha0,8'ha0,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'h80,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'h80,8'ha0,8'ha0,8'ha0,8'h80,8'ha0,8'ha0,8'ha0,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'h80,8'ha0,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'h80,8'h80,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}};

 
 	 
//////////--------------------------------------------------------------------------------------------------------------= 
always_ff@(posedge clk or negedge resetN) 
begin 
	if(!resetN) 
		RGBout <=	8'h00;  
	else begin 
		RGBout <= TRANSPARENT_ENCODING ; // default   
		if (InsideRectangle == 1'b1 && gameOver) 
			RGBout <= object_colors[offsetY][offsetX]; 		 
	end 
end 
 
//////////--------------------------------------------------------------------------------------------------------------= 
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
 
endmodule 
