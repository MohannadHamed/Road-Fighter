
 module roadFighterBitMap (

					input	logic	clk, 
					input	logic	resetN, 
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY, 
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
 
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ; 
 
 
// generating the bitmap 
 

localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel  
logic[0:63][0:127][7:0] object_colors = {
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h91,8'hb6,8'hb6,8'h91,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hf1,8'hf6,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hed,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he4,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hed,8'he0,8'he0,8'he0,8'hff,8'h71,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he4,8'hf1,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hf1,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'he0,8'he0,8'hff,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'he0,8'he0,8'he0,8'he0,8'hbf,8'h05,8'h00,8'h00,8'h6d,8'hff,8'he4,8'he0,8'he0,8'he0,8'hf6,8'hff,8'hdf,8'hdf,8'hff,8'hff,8'he4,8'he0,8'he0,8'he0,8'hfa,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hfa,8'he0,8'he0,8'he0,8'he0,8'he0,8'hed,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hf1,8'he0,8'he0,8'he0,8'he0,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h77,8'h77,8'h77,8'h77,8'h77,8'hdf,8'hed,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'hff,8'hf1,8'he0,8'he0,8'he0,8'hff,8'hff,8'h77,8'h77,8'h77,8'h77,8'hdf,8'hff,8'he0,8'he0,8'he0,8'he0,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hed,8'he0,8'he0,8'hed,8'he0,8'he0,8'he0,8'hbb,8'h2d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'hff,8'h77,8'h77,8'h77,8'h77,8'hbb,8'hff,8'hff,8'he0,8'he0,8'he0,8'hf1,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'hed,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h77,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'he0,8'he0,8'he0,8'he0,8'h9b,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hf6,8'he0,8'he0,8'he0,8'hff,8'hed,8'he0,8'he0,8'hff,8'h9b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h05,8'hf1,8'he0,8'he0,8'he0,8'hff,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'hdf,8'h77,8'h00,8'h91,8'he0,8'he0,8'he0,8'hed,8'hff,8'h77,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hf6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'hfa,8'h9b,8'hff,8'he0,8'he0,8'hed,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hf6,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h77,8'h00,8'hd6,8'he0,8'he0,8'he0,8'hf6,8'hdf,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hff,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h24,8'he0,8'he0,8'he0,8'hf1,8'hff,8'h77,8'h96,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hed,8'he0,8'he0,8'hff,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hed,8'hff,8'h77,8'h77,8'h00,8'hda,8'he0,8'he0,8'he0,8'hfb,8'hbf,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hff,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'hbb,8'h77,8'h00,8'he4,8'he0,8'he0,8'he0,8'h9b,8'h25,8'h00,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hf1,8'he0,8'he0,8'hfa,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hfa,8'hff,8'h9b,8'h77,8'h77,8'h00,8'h00,8'hfa,8'he0,8'he0,8'he0,8'hff,8'hbb,8'h05,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h6d,8'hff,8'he0,8'he0,8'he0,8'hff,8'h77,8'h05,8'h00,8'hff,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hf1,8'he0,8'he0,8'hfa,8'hbf,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'hff,8'hff,8'hff,8'he4,8'he0,8'he0,8'he0,8'hff,8'hbb,8'h77,8'h72,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hf1,8'hdf,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hfa,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'he4,8'hff,8'hff,8'hff,8'hff,8'hff,8'hf6,8'he0,8'he0,8'hf1,8'hff,8'h00,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hed,8'he0,8'he0,8'hff,8'hbb,8'h05,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h32,8'h32,8'hbb,8'hff,8'he0,8'he0,8'he0,8'hed,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h24,8'he0,8'he0,8'he0,8'he0,8'hff,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hed,8'he0,8'he0,8'he0,8'hdf,8'h77,8'h00,8'h00,8'hed,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hfa,8'h32,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'he0,8'hff,8'h05,8'h00,8'h00,8'h00,8'h00,8'he4,8'he0,8'he0,8'he0,8'hf6,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'he0,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'h6d,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hed,8'h77,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'he4,8'hff,8'h00,8'h00,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'he0,8'hff,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hff,8'he0,8'he0,8'he0,8'he0,8'hff,8'h77,8'h77,8'h00,8'hff,8'he0,8'he0,8'he0,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hf6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h24,8'hda,8'he0,8'he0,8'he0,8'hed,8'h77,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'he0,8'hdf,8'h00,8'h00,8'h00,8'h00,8'hff,8'hed,8'he0,8'he0,8'he0,8'he0,8'hfa,8'hff,8'hff,8'hfa,8'he4,8'he0,8'he0,8'he0,8'he0,8'hff,8'hbb,8'h77,8'h25,8'hff,8'hed,8'he0,8'he0,8'hff,8'hbb,8'h77,8'h77,8'h77,8'h77,8'h77,8'h77,8'h77,8'hff,8'hed,8'he0,8'he0,8'hfa,8'hdf,8'h32,8'h00,8'hda,8'he0,8'he0,8'he0,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hf1,8'he0,8'he0,8'he0,8'he0,8'hf1,8'hff,8'h77,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'he0,8'he0,8'he0,8'hf6,8'hff,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hf1,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hed,8'hff,8'h77,8'h77,8'h04,8'h00,8'hf6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'hff,8'hbb,8'h00,8'hda,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hf1,8'hbb,8'h77,8'h76,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hf1,8'he0,8'he0,8'he0,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hfa,8'hff,8'hbb,8'h77,8'h77,8'h00,8'h00,8'he4,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'he0,8'he0,8'he0,8'hf1,8'hff,8'h00,8'hda,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hff,8'hff,8'h77,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hdb,8'hdf,8'hdf,8'hdf,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hdf,8'hdf,8'hdf,8'hdf,8'h77,8'h05,8'h00,8'h00,8'h00,8'h00,8'h00,8'h9b,8'hdf,8'hff,8'hff,8'hff,8'hff,8'hff,8'hbb,8'h77,8'h77,8'h77,8'h05,8'h00,8'h00,8'h6d,8'hb6,8'hdf,8'hdf,8'hdf,8'h77,8'h77,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hdf,8'hdf,8'hdf,8'hdf,8'h32,8'h6d,8'hdb,8'hdf,8'hdf,8'hdf,8'hdf,8'hdf,8'hdf,8'hdf,8'hbf,8'hbb,8'h77,8'h77,8'h77,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h2d,8'h2d,8'h2d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h05,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h72,8'h77,8'h77,8'h76,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h2d,8'h2d,8'h2d,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h2d,8'h2d,8'h2d,8'h2d,8'h00,8'h00,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h25,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hff,8'hfa,8'hf6,8'hf1,8'hf6,8'hff,8'hff,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'h6d,8'h00,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h24,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'h00,8'h00,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'h25,8'h04,8'h00,8'hed,8'he0,8'he0,8'he0,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hfa,8'hf1,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf6,8'he0,8'he0,8'he0,8'h91,8'h04,8'hda,8'hf1,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hff,8'h2d,8'hd6,8'hf1,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hfa,8'h04,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he4,8'hf1,8'hff,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'hed,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'h00,8'h00,8'h00,8'hff,8'hed,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hff,8'hb6,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf6,8'he0,8'he0,8'he0,8'hbb,8'h77,8'hda,8'hf1,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hff,8'h9b,8'hda,8'hf1,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hba,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h77,8'h77,8'h00,8'hed,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'he0,8'hf1,8'hff,8'hff,8'hbf,8'hdf,8'hff,8'hf1,8'he0,8'he0,8'he0,8'hed,8'hff,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf6,8'he0,8'he0,8'he0,8'hbb,8'h77,8'hb6,8'hfa,8'hff,8'hff,8'hff,8'hff,8'hff,8'he0,8'he0,8'he0,8'hf1,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h77,8'hda,8'hf1,8'he0,8'he0,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdf,8'h77,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hed,8'he0,8'he0,8'he0,8'hff,8'hbf,8'h05,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'hbb,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'hed,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'he0,8'hff,8'h77,8'h77,8'h77,8'h2d,8'h2d,8'h2d,8'h96,8'hed,8'he0,8'he0,8'he0,8'hf6,8'h76,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf6,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'h00,8'h25,8'h72,8'h72,8'h72,8'h96,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h76,8'h72,8'h72,8'h72,8'h72,8'h72,8'hd6,8'hf1,8'he0,8'he0,8'hff,8'hbb,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h72,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'hff,8'h77,8'h72,8'h72,8'h72,8'h72,8'h72,8'hbb,8'hff,8'he0,8'he0,8'hed,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hed,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'h00,8'hfa,8'he0,8'he0,8'he0,8'hed,8'h9b,8'h77,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hed,8'hfb,8'hff,8'hff,8'h77,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf6,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf1,8'he0,8'he0,8'hff,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hff,8'he0,8'he0,8'hed,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hed,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'h24,8'he0,8'he0,8'he0,8'he4,8'hff,8'h77,8'h76,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h77,8'h77,8'h77,8'h77,8'h32,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf6,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf1,8'he0,8'he0,8'hff,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf1,8'he0,8'he0,8'hf6,8'hdf,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hf1,8'hf6,8'hf6,8'hf6,8'hf6,8'hf6,8'hf6,8'hf6,8'hff,8'h24,8'h00,8'h00,8'h00,8'hed,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'h91,8'he0,8'he0,8'he0,8'hf1,8'hff,8'h76,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'he0,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he0,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf1,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hf6,8'h00,8'h00,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'he0,8'he0,8'he0,8'he0,8'hff,8'h77,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hff,8'h9b,8'h00,8'h00,8'h00,8'hed,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'hd6,8'he0,8'he0,8'he0,8'hfa,8'hdf,8'h2d,8'h00,8'h00,8'h00,8'hff,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'h24,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf1,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h2d,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hf6,8'hff,8'h77,8'h77,8'h72,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hff,8'h9b,8'h00,8'h00,8'h00,8'hed,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hf6,8'hdf,8'h2d,8'h00,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'hb6,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf1,8'he0,8'he0,8'he0,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hf6,8'h77,8'h2d,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hf1,8'hfa,8'hff,8'h9b,8'h77,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'hdf,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'hbb,8'h77,8'h00,8'h00,8'h00,8'hed,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'h6d,8'he0,8'he0,8'he0,8'hed,8'hff,8'h2d,8'h00,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h77,8'h77,8'h77,8'h77,8'h77,8'h77,8'hf6,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf1,8'he0,8'he0,8'hff,8'hbb,8'h77,8'h77,8'h77,8'h77,8'h77,8'h77,8'h77,8'h77,8'h77,8'h77,8'h2d,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'hff,8'hff,8'hff,8'hff,8'he4,8'he0,8'he0,8'hf6,8'hff,8'h77,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'hbb,8'h2d,8'h05,8'h05,8'h05,8'h05,8'h05,8'h05,8'h05,8'h00,8'h00,8'h00,8'hed,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'h00,8'he4,8'he0,8'he0,8'he0,8'hff,8'h72,8'h00,8'h00,8'h00,8'h00,8'h25,8'h77,8'h77,8'hff,8'hf1,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf6,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf1,8'he0,8'he0,8'hff,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'hff,8'h77,8'h32,8'h32,8'hbb,8'he0,8'he0,8'he0,8'he0,8'hff,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hed,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'h00,8'hff,8'he0,8'he0,8'he0,8'he0,8'hdf,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hf1,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf6,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf1,8'he0,8'he0,8'hff,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'hff,8'hed,8'he0,8'he0,8'he0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hed,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'h00,8'hff,8'hf1,8'he0,8'he0,8'he0,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hff,8'hed,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf6,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf1,8'he0,8'he0,8'hff,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h6d,8'hff,8'he0,8'he0,8'he0,8'he4,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hed,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'h00,8'h00,8'hb1,8'he0,8'he0,8'he0,8'he0,8'he0,8'hfa,8'hff,8'hff,8'hff,8'hf1,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf6,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf1,8'he0,8'he0,8'hfa,8'hfb,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hfa,8'hff,8'h24,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'hfb,8'hdf,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hed,8'he0,8'he0,8'he0,8'h9b,8'h77,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'he4,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hf1,8'hff,8'hff,8'h77,8'h77,8'h00,8'hb6,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf6,8'he0,8'he0,8'he0,8'hbb,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'he0,8'he0,8'he0,8'hf1,8'h77,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf1,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'he0,8'hff,8'h9b,8'h00,8'h00,8'hf1,8'he0,8'he0,8'he0,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hfa,8'he0,8'he0,8'he0,8'hf6,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'hf6,8'hf6,8'hf6,8'hff,8'hbb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hf6,8'hf6,8'hf6,8'h9b,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h72,8'hff,8'hff,8'hf1,8'hed,8'he0,8'he4,8'hed,8'hf6,8'hff,8'hff,8'h77,8'h77,8'h77,8'h2d,8'h00,8'h00,8'hb6,8'hf6,8'hf6,8'hf6,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hf6,8'hf6,8'hf6,8'hbb,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hf6,8'hf6,8'hf6,8'hfa,8'h77,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hfa,8'hf6,8'hf6,8'hf6,8'hf6,8'hf6,8'hf6,8'hf6,8'hf6,8'hf6,8'hf6,8'hf6,8'hf6,8'hf6,8'hff,8'h9b,8'h00,8'h00,8'hfa,8'hf6,8'hf6,8'hf6,8'hff,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hf6,8'hf6,8'hf6,8'hf6,8'hfa,8'h76,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h6d,8'hdb,8'hdf,8'hdf,8'hdf,8'h9b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hdf,8'hdf,8'hdf,8'h77,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h77,8'hbb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hdf,8'h77,8'h77,8'h77,8'h77,8'h72,8'h00,8'h00,8'h00,8'h6d,8'hdb,8'hdf,8'hdf,8'hdf,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hdb,8'hdf,8'hdf,8'h9b,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hdf,8'hdf,8'hdf,8'h77,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hb6,8'hdf,8'hdf,8'hdf,8'hdf,8'hdf,8'hdf,8'hdf,8'hdf,8'hdf,8'hdf,8'hdf,8'hdf,8'hdf,8'hdf,8'h77,8'h00,8'h00,8'hb6,8'hdb,8'hdf,8'hdf,8'hdf,8'h77,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdf,8'hdf,8'hdf,8'hdf,8'hdf,8'h77,8'h05,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h2d,8'h2d,8'h2d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h05,8'h2d,8'h2d,8'h2d,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h05,8'h2d,8'h76,8'h77,8'h77,8'h76,8'h2d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h2d,8'h2d,8'h2d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h2d,8'h2d,8'h2d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h2d,8'h2d,8'h2d,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h2d,8'h2d,8'h2d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h05,8'h2d,8'h2d,8'h2d,8'h2d,8'h2d,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}};

 
 	 
//////////--------------------------------------------------------------------------------------------------------------= 
always_ff@(posedge clk or negedge resetN) 
begin 
	if(!resetN) begin 
		RGBout <=	8'h00; 
	end 
	else begin 
		RGBout <= TRANSPARENT_ENCODING ; // default   
		if (InsideRectangle == 1'b1 ) 
			RGBout <= object_colors[offsetY][offsetX]; 
		 
	end 
end 
 
//////////--------------------------------------------------------------------------------------------------------------= 
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
 
endmodule 
